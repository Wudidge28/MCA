BZh91AY&SY�RV �߀Ryg����������P޸ʎ�;X �DhBmS�I�F����  5=@m@�2�S�zF�F��@i��@ $D�#"=#��F��Pz� ��dɡ��рFa `&�4��$�F�� (jzO
~�z���4P24ڗ�$̆8�g�	�(�Ji%�Q/oÜC�=DAS���7��j.�ʥ�&�\�v�	���̣0���+dJ����V����r�d`W,��Ս���Y�:z���i�f�d�OfI�;��%l����~ao��w��%	� W6�ǁJ�0�7	��٩�yn�;�ؘȄ�@��I##G���BE���S�U���ZY���w@�ؘUH�ss[󫆈
��*Pj��54����
�L�ʞ(��e��=�k�S��i{%}��(!��$��}K�����Cl�6��y$p[�A��e��)D��`��4���A��Zi�� T��X�S�ߒQ���b���\&w3R"Q��AΪ.^��`�#	#O4�m45��ͭ]����P&�{<QO��]

�q@�73,1�T�Az�S�)&����w��'G 7H�O�^ v"U	u��@;O��M��p�U�]�z�''>�D��a��1�n��~����Ƶ��#@5/�sf�1�80!+rٺ�mF��Q;�,���Z&4Lq��?I@��Z̖��ʌBt��E�h1���D�h�!D(�,\ș���S1Ņ�����mg"v��Q��	�xY=y�J	|Y6�TaO��G�z �8:����C/9!iC�=���!�fV<Nq��8ɂb��
ך\�}=\2�K�L��h/2G��v-��Pc�Bdo�m�&��:�kf��;(n��O,XC����Ǖ!��3�TriK�Y2�Ҹ��9�$Y�6@�L�&jIF�x�m�Z�cJD�߉���ɞ��J�q�q6�O��*(�P�3�P��=rE��&ī��j&&�i;f���e���H��#��fp.��-�<�����g�b��H%~��\�u�j�Q�
�35�{����#�iw�z<���2ֹ�(d�8@c��$Q�����}��Q*EHŀ��c$�����. l�\�0x#Ea�*%�h��
�`f&YĿ�[*��Vظ�ڡ��ƨF��q͚�C+����:<�h6����gEy�qyz��"����)*�`̋hm�zђiP8��ȱ��.�p� =���